// neccesary parameters for verilog modules 
`define N_CHANNEL_EN 32
